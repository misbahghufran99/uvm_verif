 interface new_cuboid_inp_intf (input clk);

  logic [16-1:0] in_data;
  logic          valid ;
  logic          start ;

endinterface
