 interface new_cuboid_out_intf (input clk);

  logic [32-1:0]  out_data ;
  logic          valid;
  logic           start;

endinterface